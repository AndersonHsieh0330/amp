** sch_path: /home/andersonhsieh/repos/projects/amp/characterization/characterization.sch
**.subckt characterization
XM3 GND net1 net2 net2 sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
Vgs net1 GND 1.8
Vds_p net2 GND 0.9
**** begin user architecture code

.control
    save all
    +@m.xm1.msky130_fd_pr__nfet_01v8[id] @m.xm1.msky130_fd_pr__nfet_01v8[gm]
    +@m.xm2.msky130_fd_pr__pfet_01v8[id] @m.xm2.msky130_fd_pr__pfet_01v8[gm]
    dc Vgs 0 2 0.1
    write out.raw
.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
